module bcdadder(a,b,cou,sum);
    input[3:0] a,b;
    output[3:0] sum;
    output cou;
    always @(*)
      if(sum > 4'd9)
        
        
    
    
endmodule



